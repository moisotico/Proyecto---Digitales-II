`timescale 1ns/1ps

module gen_clk(
	clk_8f, rst, enb
	clk_2f, clk_f	
);




endmodule
